Divisor_CLK_inst : Divisor_CLK PORT MAP (
		clock	 => clock_sig,
		cout	 => cout_sig,
		q	 => q_sig
	);
