CLOCK_MINUTOS_inst : CLOCK_MINUTOS PORT MAP (
		clock	 => clock_sig,
		cout	 => cout_sig,
		q	 => q_sig
	);
